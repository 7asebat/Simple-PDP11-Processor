Library ieee;
Use ieee.std_logic_1164.all;
use ieee.numeric_std.ALL;
use IEEE.math_real.all;

ENTITY nmROM IS 
	PORT(
    address: IN std_logic_vector(integer(ceil(log2(real(65536))))-1 DOWNTO 0);
    dataOut: OUT std_logic_vector(21-1 DOWNTO 0)
  ); 
END ENTITY;

ARCHITECTURE main OF nmRom IS
  CONSTANT n: integer := 256; -- ROM size
  CONSTANT m: integer := 21; -- Control Signal Width
  TYPE rom_type IS ARRAY(0 TO n-1) of std_logic_vector(m-1 DOWNTO 0);
  SIGNAL rom: rom_type := (
    0 => "000101101000001011100",
    1 => "001100100001111000010",
    2 => "001001000001111000000",
    3 => "000000000001111000001",
    4 => "010000000101111000000",
    5 => "000000000001111000001",
    6 => "010000001001111010010",
    7 => "000000000001111000001",
    8 => "010001101000001001110",
    9 => "001110000001111000010",
    10 => "000000000001111000001",
    11 => "010001100000010001100",
    12 => "001110001001111010010",
    13 => "000000000001111000001",
    14 => "000101101000001011100",
    15 => "001100100001111000010",
    16 => "001000000011111000000",
    17 => "010001100000001000000",
    18 => "001100001001111010010",
    19 => "000000000001111000001",
    20 => "001000001001111010010",
    21 => "001000000101111000000",
    22 => "000000000001111000001",
    23 => "010100000111111000000",
    24 => "000000000001111000001",
    25 => "010100001001111010010",
    26 => "000000000001111000001",
    27 => "010101101000001011100",
    28 => "001110100001111000010",
    29 => "000000000001111000001",
    30 => "010101100000010001100",
    31 => "001110101001111010010",
    32 => "000000000001111000001",
    33 => "000101101000001011100",
    34 => "001100100001111000010",
    35 => "001000000011111000000",
    36 => "010101100000001000000",
    37 => "001100001001111010010",
    38 => "000000000001111000001",
    39 => "001000001001111010010",
    40 => "001000000111111000000",
    41 => "000000000001111000001",
    42 => "011001100000001001000",
    43 => "000000000001111000001",
    44 => "011000000011111000000",
    45 => "011101100000001000000",
    46 => "000000000001111000001",
    47 => "011000000011111000000",
    48 => "011101100000001000100",
    49 => "000000000001111000001",
    50 => "011000000011111000000",
    51 => "011101100000010000100",
    52 => "000000000001111000001",
    53 => "011000000011111000000",
    54 => "011101100000010000000",
    55 => "000000000001111000001",
    56 => "011000000011111000000",
    57 => "011101100000100000000",
    58 => "000000000001111000001",
    59 => "011000000011111000000",
    60 => "011101100000101000000",
    61 => "000000000001111000001",
    62 => "011000000011111000000",
    63 => "011101100000110000000",
    64 => "000000000001111000001",
    65 => "011000000011111000000",
    66 => "011101100000010000000",
    67 => "000000000001111000001",
    68 => "011101100000001001100",
    69 => "000000000001111000001",
    70 => "011101100000010001100",
    71 => "000000000001111000001",
    72 => "011101100000100001000",
    73 => "000000000001111000001",
    74 => "011101100000111000000",
    75 => "000000000001111000001",
    76 => "011101100001000000000",
    77 => "000000000001111000001",
    78 => "011101100001001000000",
    79 => "000000000001111000001",
    80 => "011101100001011000000",
    81 => "000000000001111000001",
    82 => "011101100001100000000",
    83 => "000000000001111000001",
    84 => "011101100001101000000",
    85 => "000000000001111000001",
    86 => "100000000101111000000",
    87 => "000100000111111000000",
    88 => "000000000001111000001",
    89 => "001100100001111000000",
    90 => "000000000001111000001",
    91 => "000000000000000000000",
    92 => "000000000000000000000",
    93 => "000000000001111000001",
    94 => "000101101000001011100",
    95 => "001100100001111000010",
    96 => "001000000101111000010",
    97 => "000100010001111000000",
    98 => "000000000001111000001",
    99 => "100000100001111000000",
    100 => "000000000001111000001",
    101 => "100100010001111000000",
    102 => "000000000001111000001",
    103 => "000100010001111000000",
    104 => "101001100000010001100",
    105 => "001111101001111100010",
    106 => "101100100001111000000",
    107 => "000000000001111000001",
    108 => "101001101000001011100",
    109 => "001111100001111000010",
    110 => "001000100001111000000",
    111 => "000000000001111000001",
    112 => "101001101000001011100",
    113 => "001111100001111000010",
    114 => "001011000001111000000",
    115 => "000000000001111000001",
    116 => "101001100000010001100",
    117 => "001111101001111100010",
    118 => "000000000001111000001",
    119 => "001110100001111000000",
    120 => "000000000001111000001",
    121 => "001100010001111100010",
    122 => "000000000001111000001",
    OTHERS => ("000000000000000000000")
  );
BEGIN
  dataOut <= rom(to_integer(unsigned(address)));
END ARCHITECTURE;