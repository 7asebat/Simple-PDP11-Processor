Library ieee;
Use ieee.std_logic_1164.all;
use ieee.numeric_std.ALL;
use IEEE.math_real.all;

ENTITY nmROM IS 
	PORT(
    address: IN std_logic_vector(integer(ceil(log2(real(n))))-1 DOWNTO 0);
    dataOut: OUT std_logic_vector(m-1 DOWNTO 0)
  ); 
END ENTITY;

ARCHITECTURE main OF nmRam IS
  CONSTANT n: integer := 128; -- ROM size
  CONSTANT m: integer := 21; -- Control Signal Width
  TYPE rom_type IS ARRAY(0 TO n-1) of std_logic_vector(m-1 DOWNTO 0);
  SIGNAL rom: rom_type := (
    0 => "000101101000001011100",
    1 => "001100100000000000010",
    2 => "001001000000000000000",
    3 => "000000000000000000001",
    4 => "010000000100000000000",
    5 => "000000000000000000001",
    6 => "010000001000000010010",
    7 => "000000000000000000001",
    8 => "010001101000001001110",
    9 => "001110000000000000000",
    10 => "000000000000000000001",
    11 => "010001100000010001100",
    12 => "001110001000000010010",
    13 => "000000000000000000001",
    14 => "000101101000001011100",
    15 => "001100100000000000000",
    16 => "001000000010000000000",
    17 => "010001100000001000000",
    18 => "001100001000000010010",
    19 => "000000000000000000001",
    20 => "001000001000000010010",
    21 => "001000000100000000000",
    22 => "000000000000000000001",
    23 => "010100000110000000000",
    24 => "000000000000000000001",
    25 => "010100001000000010010",
    26 => "000000000000000000001",
    27 => "010101101000001011100",
    28 => "001110100000000000010",
    29 => "000000000000000000001",
    30 => "010101100000010001100",
    31 => "001110101000000010010",
    32 => "000000000000000000001",
    33 => "000101101000001011100",
    34 => "001100100000000000010",
    35 => "001000000010000000000",
    36 => "010101100000001000000",
    37 => "001100001000000010010",
    38 => "000000000000000000001",
    39 => "001000001000000010010",
    40 => "001000000110000000000",
    41 => "000000000000000000001",
    42 => "011011000110000000000",
    43 => "000000000000000000001",
    44 => "011000000010000000000",
    45 => "011101100000001000000",
    46 => "000000000000000000001",
    47 => "011000000010000000000",
    48 => "011101100000001000100",
    49 => "000000000000000000001",
    50 => "011000000010000000000",
    51 => "011101100000010000100",
    52 => "000000000000000000001",
    53 => "011000000010000000000",
    54 => "011101100000010000000",
    55 => "000000000000000000001",
    56 => "011000000010000000000",
    57 => "011101100000100000000",
    58 => "000000000000000000001",
    59 => "011000000010000000000",
    60 => "011101100000101000000",
    61 => "000000000000000000001",
    62 => "011000000010000000000",
    63 => "011101100000110000000",
    64 => "000000000000000000001",
    65 => "011000000010000000000",
    66 => "011101100000010000000",
    67 => "000000000000000000001",
    68 => "011101100000001001100",
    69 => "000000000000000000001",
    70 => "011101100000010001100",
    71 => "000000000000000000001",
    72 => "011101100000100001000",
    73 => "000000000000000000001",
    74 => "011101100000111000000",
    75 => "000000000000000000001",
    76 => "011101100001000000000",
    77 => "000000000000000000001",
    78 => "011101100001001000000",
    79 => "000000000000000000001",
    80 => "011101100001011000000",
    81 => "000000000000000000001",
    82 => "011101100001100000000",
    83 => "000000000000000000001",
    84 => "011101100001101000000",
    85 => "000000000000000000001",
    86 => "100000000100000000000",
    87 => "000100000110000000000",
    88 => "000000000000000000001",
    89 => "001100100000000000000",
    90 => "000000000000000000001",
    91 => "000000000000000000001",
    92 => "000101101000001011100",
    93 => "001100100000000000010",
    94 => "001000000100000000010",
    95 => "000100010000000000000",
    96 => "000000000000000000001",
    97 => "100000100000000000000",
    98 => "000000000000000000001",
    99 => "100100010000000000000",
    100 => "000000000000000000001",
    101 => "000100010000000000000",
    102 => "101001100000010001100",
    103 => "001111101000000100010",
    104 => "101100100000000000000",
    105 => "000000000000000000001",
    106 => "101001101000001011110",
    107 => "001111100000000000000",
    108 => "001000100000000000000",
    109 => "000000000000000000001",
    110 => "101001101000001011100",
    111 => "001111100000000000010",
    112 => "001011000000000000000",
    113 => "000000000000000000001",
    114 => "101001100000010001100",
    115 => "001111101000000100010",
    116 => "000000000000000000001",
    117 => "001110100000000000000",
    118 => "000000000000000000001",
    119 => "001100010000000100010",
    120 => "000000000000000000001",
  );
BEGIN
  dataOut <= rom(to_integer(unsigned(address)));
END ARCHITECTURE;