Library ieee;
Use ieee.std_logic_1164.all;
use ieee.numeric_std.ALL;
use IEEE.math_real.all;

ENTITY nmROM IS 
	PORT(
    address: IN std_logic_vector(integer(ceil(log2(real(n))))-1 DOWNTO 0);
    dataOut: OUT std_logic_vector(m-1 DOWNTO 0)
  ); 
END ENTITY;

ARCHITECTURE main OF nmRam IS
  CONSTANT n: integer := 128; -- ROM size
  CONSTANT m: integer := 21; -- Control Signal Width
  TYPE rom_type IS ARRAY(0 TO n-1) of std_logic_vector(m-1 DOWNTO 0);
  SIGNAL rom: rom_type := (
    0 => "000101101000001011100",
    1 => "001100100000000000010",
    2 => "001001000000000000000",
    3 => "000000000000000000001",
    4 => "010000000100000000000",
    5 => "000000000000000000001",
    6 => "010000001000000010010",
    7 => "000000000000000000001",
    8 => "010001101000001001110",
    9 => "001110000000000000000",
    10 => "000000000000000000001",
    11 => "010001100000010001100",
    12 => "001110001000000010010",
    13 => "000000000000000000001",
    14 => "000101101000001011100",
    15 => "001100100000000000000",
    16 => "001000000010000000000",
    17 => "010001100000001000000",
    18 => "001100001000000010010",
    19 => "000000000000000000001",
    20 => "001000001000000010010",
    21 => "001000000100000000000",
    22 => "010100000110000000000",
    23 => "000000000000000000001",
    24 => "010100001000000010010",
    25 => "000000000000000000001",
    26 => "010101101000001011100",
    27 => "001110100000000000010",
    28 => "000000000000000000001",
    29 => "010101100000010001100",
    30 => "001110101000000010010",
    31 => "000000000000000000001",
    32 => "000101101000001011100",
    33 => "001100100000000000010",
    34 => "001000000010000000000",
    35 => "010101100000001000000",
    36 => "001100001000000010010",
    37 => "000000000000000000001",
    38 => "001000001000000010010",
    39 => "001000000110000000000",
    40 => "000000000000000000001",
    41 => "011011000110000000000",
    42 => "000000000000000000001",
    43 => "011000000010000000000",
    44 => "011101100000001000000",
    45 => "000000000000000000001",
    46 => "011000000010000000000",
    47 => "011101100000001000100",
    48 => "000000000000000000001",
    49 => "011000000010000000000",
    50 => "011101100000010000100",
    51 => "000000000000000000001",
    52 => "011000000010000000000",
    53 => "011101100000010000000",
    54 => "000000000000000000001",
    55 => "011000000010000000000",
    56 => "011101100000100000000",
    57 => "000000000000000000001",
    58 => "011000000010000000000",
    59 => "011101100000101000000",
    60 => "000000000000000000001",
    61 => "011000000010000000000",
    62 => "011101100000110000000",
    63 => "000000000000000000001",
    64 => "011000000010000000000",
    65 => "011101100000010000000",
    66 => "000000000000000000001",
    67 => "011101100000001001100",
    68 => "000000000000000000001",
    69 => "011101100000010001100",
    70 => "000000000000000000001",
    71 => "011101100000100001000",
    72 => "000000000000000000001",
    73 => "011101100000111000000",
    74 => "000000000000000000001",
    75 => "011101100001000000000",
    76 => "000000000000000000001",
    77 => "011101100001001000000",
    78 => "000000000000000000001",
    79 => "011101100001011000000",
    80 => "000000000000000000001",
    81 => "011101100001100000000",
    82 => "000000000000000000001",
    83 => "011101100001101000000",
    84 => "000000000000000000001",
    85 => "100000000100000000000",
    86 => "000100000110000000000",
    87 => "000000000000000000001",
    88 => "001100100000000000000",
    89 => "000000000000000000001",
    90 => "000000000000000000001",
    91 => "000101101000001011100",
    92 => "001100100000000000010",
    93 => "001000000100000000010",
    94 => "000100010000000000000",
    95 => "000000000000000000001",
    96 => "100000100000000000000",
    97 => "000000000000000000001",
    98 => "100100010000000000000",
    99 => "000000000000000000001",
    100 => "000100010000000000000",
    101 => "101001100000010001100",
    102 => "001111101000000100010",
    103 => "101100100000000000000",
    104 => "000000000000000000001",
    105 => "101001101000001011110",
    106 => "001111100000000000000",
    107 => "001000100000000000000",
    108 => "000000000000000000001",
    109 => "101001101000001011100",
    110 => "001111100000000000010",
    111 => "001011000000000000000",
    112 => "000000000000000000001",
    113 => "101001100000010001100",
    114 => "001111101000000100010",
    115 => "000000000000000000001",
    116 => "001110100000000000000",
    117 => "000000000000000000001",
    118 => "001100010000000100010",
    119 => "000000000000000000001",
  );
BEGIN
  dataOut <= rom(to_integer(unsigned(address)));
END ARCHITECTURE;