-- Working processor here
