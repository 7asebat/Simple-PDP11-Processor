Library ieee;
Use ieee.std_logic_1164.all;
use ieee.numeric_std.ALL;
use IEEE.math_real.all;

ENTITY nmRam IS 
  GENERIC(
    n: INTEGER := 32;
    m: INTEGER := 32
  );
  PORT(
    clk: IN std_logic;
    MFC: OUT std_logic;
    read: in std_logic;
    write: in std_logic;
    address: IN std_logic_vector(integer(ceil(log2(real(n))))-1 DOWNTO 0);
    dataIn: IN std_logic_vector(m-1 DOWNTO 0);
    dataOut: OUT std_logic_vector(m-1 DOWNTO 0)
  ); 
END ENTITY;

ARCHITECTURE main OF nmRam IS
  constant DELAY: integer := 2;

  TYPE ram_type IS ARRAY(0 TO n-1) of std_logic_vector(m-1 DOWNTO 0);
  SIGNAL ram: ram_type := (
    -- initialize here 
    0 => ("0000010111000000"),
    1 => ("0000000000000001"),
    2 => ("1100000000000010"),
    3 => ("0000010111000000"),
    4 => ("0000000000000010"),
    5 => ("0000010111000000"),
    6 => ("0000000000000011"),
    7 => ("1001001000000100"),
    8 => ("1100100000000010"),
    9 => ("0000010111000000"),
    10 => ("0000000000000100"),
    11 => ("0000010111000000"),
    12 => ("0000000000000101"),
    13 => ("0001010111000001"),
    14 => ("0000000000000001"),
    15 => ("1101000000000010"),
    16 => ("0000010111000000"),
    17 => ("0000000000000110"),
    18 => ("0000010111000000"),
    19 => ("0000000000000111"),
    20 => ("0000010111000001"),
    21 => ("0000000000000101"),
    22 => ("0000010111000010"),
    23 => ("0000000000000110"),
    24 => ("1000000001000010"),
    25 => ("1101100000000010"),
    26 => ("0000010111000000"),
    27 => ("0000000000001000"),
    28 => ("0000010111000000"),
    29 => ("0000000000001001"),
    30 => ("0000010111000001"),
    31 => ("0000000000000110"),
    32 => ("0000010111000010"),
    33 => ("0000000000000110"),
    34 => ("1000000001000010"),
    35 => ("1110000000000010"),
    36 => ("0000010111000000"),
    37 => ("0000000000001010"),
    38 => ("0000010111000000"),
    39 => ("0000000000001011"),
    40 => ("0000010111000001"),
    41 => ("0000000000000101"),
    42 => ("0000010111000010"),
    43 => ("0000000000000110"),
    44 => ("1000000001000010"),
    45 => ("1110000000000010"),
    46 => ("0000010111000000"),
    47 => ("0000000000001100"),
    48 => ("0000010111000000"),
    49 => ("0000000000001101"),
    50 => ("0000010111000001"),
    51 => ("0000000000000111"),
    52 => ("0000010111000010"),
    53 => ("0000000000000110"),
    54 => ("1000000001000010"),
    55 => ("1110100000000010"),
    56 => ("0000010111000000"),
    57 => ("0000000000001110"),
    58 => ("0000010111000000"),
    59 => ("0000000000001111"),
    60 => ("0000010111000001"),
    61 => ("0000000000000111"),
    62 => ("0000010111000010"),
    63 => ("0000000000000110"),
    64 => ("1000000001000010"),
    65 => ("1111000000000010"),
    66 => ("0000010111000000"),
    67 => ("0000000000010000"),
    68 => ("0000010111000000"),
    69 => ("0000000000010001"),
    70 => ("0000010111000001"),
    71 => ("0000000000000110"),
    72 => ("0000010111000010"),
    73 => ("0000000000000110"),
    74 => ("1000000001000010"),
    75 => ("1111000000000010"),
    76 => ("0000010111000000"),
    77 => ("0000000000010010"),
    78 => ("0000010111000000"),
    79 => ("0000000000010011"),
    80 => ("1010000000000000"),
    OTHERS => ((m-1 DOWNTO 8 => '0') & X"00")
  );
  SIGNAL s_mfc: std_logic := '0';
BEGIN

MFC <= s_mfc;

-- Delay write operation by two clock cycles
PROCESS(clk, read, write)
  variable v_delay: natural range 0 to DELAY := 0;
BEGIN
  IF(read = '0' AND write = '0') THEN
    v_delay := 0;
  END IF;

  IF(rising_edge(clk)) THEN
    v_delay := v_delay + 1;
    
    if v_delay = DELAY then
      v_delay := 0;

      if write = '1' then
        ram(to_integer(unsigned(address))) <= dataIn;
        dataOut <= dataIn;
      elsif read = '1' then
        dataOut <= ram(to_integer(unsigned(address)));
      end if;

      s_mfc <= '1';
    else
      s_mfc <= '0';
    end if;
  end if;

end process;
end architecture;